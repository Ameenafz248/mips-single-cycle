module tb;
reg clk;
reg reset;
wire [63:0] writedata, dataadr;
wire memwrite;
// instantiate device to be tested
top dut(clk, reset, writedata, dataadr, memwrite);
// initialize test
// initial begin
//     $monitor("instr: %h", instr);
// end
initial
begin
reset <= 1; # 22; reset <= 0;
end
// generate clock to sequence tests
always
begin
clk <= 1; # 5; clk <= 0; # 5;
end
// check results
always @ (negedge clk)begin
if (memwrite) begin
if (dataadr === 20 && writedata === 1000) begin
$display ("Simulation succeeded");
$stop;
end else if (dataadr !== 80) begin
$display ("Failed hehe %h and %h",writedata,dataadr);
$finish;
end
end
end
endmodule